----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 15.06.2022 09:56:09
-- Design Name: 
-- Module Name: tb_mov_avg_filter - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity tb_mov_avg_filter is
--  Port ( );
end tb_mov_avg_filter;

architecture Behavioral of tb_mov_avg_filter is
component mov_avg_filter is
    generic(M: integer := 8);
    Port (clk: in std_logic; input: in std_logic_vector(15 downto 0); output: out std_logic_vector(15 downto 0) );
end component;
type sample_array is array(0 to 255) of signed(15 downto 0); 
signal samples: sample_array := (
"0000011100101100",
"0011001110010010",
"0010000110001011",
"0100010010110100",
"0101001100011011",
"0100111101010110",
"0110110111010100",
"0101000101110011",
"0110111011010110",
"0110111011000111",
"0110101001101100",
"1000011000010011",
"0111011001000000",
"0111101111000000",
"1001101101010110",
"0111111101100001",
"1001001100011110",
"0111111101100001",
"0111110110001001",
"1001101011010101",
"1000101101011101",
"0111000011100001",
"0111001001010100",
"0110011010101000",
"0101110011101111",
"0110101001100101",
"0101001110010000",
"0101001100110111",
"0011100000000100",
"0011011000011101",
"0010101000100110",
"0010011001100000",
"0000011001011000",
"0000011010011110",
"0000000110111100",
"1110011111111110",
"1101111011001111",
"1101111101011000",
"1101110011111001",
"1101010010100100",
"1010101111000001",
"1011000001011011",
"1001010110111011",
"1011010100100011",
"1001010110010110",
"1010011110110101",
"1010001000001000",
"1001111100001000",
"1001100100100001",
"1001001100001001",
"1001111101101000",
"1001111001101101",
"1000111010010000",
"1010101001111011",
"1011000111011100",
"1011001101101000",
"1011000100000111",
"1010111101001011",
"1101110110101101",
"1100011111101101",
"1101011100110100",
"1110110101000110",
"0000000010110110",
"0000011010101001",
"0000010001101111",
"0001011001110010",
"0011110111111011",
"0011111111000101",
"0100001000000010",
"0011111000100110",
"0100110110100100",
"0110010010001001",
"0101110101011010",
"0111110000110000",
"0111001101001111",
"1000001111110111",
"0111011001000000",
"1001001011001110",
"1000001110100101",
"0111111101100001",
"0111111111111111",
"0111111101100001",
"0111110110001001",
"0111101001111100",
"0111111001000110",
"1000111110100001",
"0111001000011010",
"0110110010100101",
"0101101011011110",
"0111001001001010",
"0101010000111001",
"0100101001011011",
"0100010000000010",
"0011000001011111",
"0010111101111100",
"0010100010110110",
"0001111011110000",
"1111010001010110",
"1111001111001000",
"1111100110001111",
"1101011100001010",
"1110001011110000",
"1101001111000110",
"1100001111111010",
"1011101000111010",
"1100000001011110",
"1010000011100010",
"1010011100001000",
"1010010001100110",
"1010101111111011",
"1000001100000100",
"1000111101110110",
"1000100101000011",
"1001011110001101",
"1000011001010011",
"1010010011001110",
"1001100100111110",
"1001100011000111",
"1010100110011111",
"1010001111110110",
"1100100100011010",
"1011110111111010",
"1011101010100011",
"1101011110000010",
"1110000110110110",
"1110010001000000",
"0000101111111000",
"0001001100101111",
"0010000111101011",
"0000110010010010",
"0011011100110011",
"0100011001010110",
"0011001001010001",
"0011110100000110",
"0110101100011101",
"0101000100110011",
"0101110011010111",
"0110001011110001",
"1000000000000011",
"1000010010011101",
"0111011001000000",
"0111101001111100",
"0111110110001001",
"0111111101100001",
"1001110011110001",
"1000111011110100",
"0111110110001001",
"1000001011000111",
"0111011001000000",
"0111010101100110",
"0110101001101100",
"0110001011110001",
"0101101010000001",
"0101000100110011",
"0110001001011011",
"0100011010000001",
"0011110000111001",
"0010011101000010",
"0001111011101010",
"0001100010111100",
"0000111010100000",
"1111101100111111",
"0000100101111101",
"1111101010110001",
"1110000000001110",
"1101100100111001",
"1100100000001011",
"1101001110010001",
"1100010110111011",
"1010011110100001",
"1001110011110010",
"1001100010101110",
"1001100011111111",
"1001111000110010",
"1000111110101001",
"1001111101100101",
"1000101111101110",
"1010000011110011",
"1001010001010110",
"1010010000010000",
"1001010111000100",
"1001110010000101",
"1011001001001011",
"1010011100000110",
"1100101100010110",
"1010111110011001",
"1011110101100001",
"1101111001001000",
"1110111101010010",
"1110111110101100",
"1111011001010011",
"0000001101010110",
"0000101000010000",
"0001011100000100",
"0001101011110101",
"0010101101011000",
"0011110000101010",
"0101010010001000",
"0101000010110000",
"0101000100110011",
"0110000110101101",
"0110001011110001",
"0110111011100000",
"0111000011100001",
"0111011001000000",
"0111101001111100",
"0111110110001001",
"0111111101100001",
"1000010110010001",
"1000000111110010",
"0111110110001001",
"1001001101001010",
"0111011001000000",
"1001011010001100",
"0110101001101100",
"0110111101100011",
"0110010100010101",
"0110010011111001",
"0100111100000110",
"0100100001001000",
"0011100011001001",
"0011010011000110",
"0011000010010010",
"0010010110100100",
"0001110000011010",
"1111010101011001",
"0000100100011011",
"1111000000110100",
"1101100101111100",
"1100011010010011",
"1011100101101010",
"1100100000111001",
"1010011001100110",
"1001111110110101",
"1011001111101011",
"1010101100100101",
"1000101110000001",
"1000110110001010",
"1000101011100111",
"1001001110100101",
"1000111011100010",
"1001010000001001",
"1001101010000010",
"1001011000110011",
"1001000101110011",
"1011001101110011",
"1001100110100000",
"1011100111100110",
"1010111110001011",
"1011011100011010",
"1101011101101001",
"1101011000111111",
"1110011001000110",
"1111011110101000",
"0000001010110111",
"1111101101111110"

);
signal clk: std_logic := '1';
constant cycles: integer := 256;
constant T: time := 20 ns;
signal input: std_logic_vector(15 downto 0) := (others => '0');
signal output: std_logic_vector(15 downto 0) := (others => '0');
begin
tb: mov_avg_filter port map(clk => clk, input => input, output => output);
process
begin
    for i in 0 to cycles - 1 loop
      clk <= '0';
      wait for T / 2;
      clk <= '1';
      wait for T / 2;
    end loop;
    wait;
    
end process;


process(clk)
variable i: integer := 0;
begin
    if rising_edge(clk) then
        input <= std_logic_vector(samples(i));
        i := i + 1;
    end if;
end process;


end Behavioral;
